library verilog;
use verilog.vl_types.all;
entity celula_vlg_vec_tst is
end celula_vlg_vec_tst;
