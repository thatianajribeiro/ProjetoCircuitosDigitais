library verilog;
use verilog.vl_types.all;
entity soma_vlg_vec_tst is
end soma_vlg_vec_tst;
