    library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity decodificador is
    Port ( instrucao : in  STD_LOGIC_VECTOR (7 downto 0);
    	   out_decod : out STD_LOGIC_VECTOR(10 downto 0));
end decodificador;

architecture archdecodificador of decodificador is

begin	
	process (instrucao)
	begin
		-- Inicializa todos em 0
		out_decod <= "00000000000";
		case instrucao(7 downto 4) is
			when "0000" => out_decod <= "10000000000"; --nop;
			when "0001" => out_decod <= "01000000000"; --sta;
			when "0010" => out_decod <= "00100000000"; --lda;
			when "0011" => out_decod <= "00010000000"; --add;
			when "0100" => out_decod <= "00001000000"; --or;
			when "0101" => out_decod <= "00000100000"; --and;
			when "0110" => out_decod <= "00000010000"; --not;
			when "1000" => out_decod <= "00000001000"; --jmp;
			when "1001" => out_decod <= "00000000100"; --jn;
			when "1010" => out_decod <= "00000000010"; --jz;
			when "1111" => out_decod <= "00000000001"; --hlt <= '1';
			when others => out_decod <= "00000000000"; 
		end case;
	end process;
end archdecodificador;